magic
tech sky130A
timestamp 1687720305
<< nwell >>
rect -315 180 90 320
<< nmos >>
rect -195 25 -180 125
rect 5 25 20 125
<< pmos >>
rect -195 200 -180 300
rect 5 200 20 300
<< ndiff >>
rect -245 105 -195 125
rect -245 45 -230 105
rect -210 45 -195 105
rect -245 25 -195 45
rect -180 105 -130 125
rect -180 45 -165 105
rect -145 45 -130 105
rect -180 25 -130 45
rect -45 105 5 125
rect -45 45 -30 105
rect -10 45 5 105
rect -45 25 5 45
rect 20 105 70 125
rect 20 45 35 105
rect 55 45 70 105
rect 20 25 70 45
<< pdiff >>
rect -245 280 -195 300
rect -245 220 -230 280
rect -210 220 -195 280
rect -245 200 -195 220
rect -180 280 -130 300
rect -180 220 -165 280
rect -145 220 -130 280
rect -180 200 -130 220
rect -45 280 5 300
rect -45 220 -30 280
rect -10 220 5 280
rect -45 200 5 220
rect 20 280 70 300
rect 20 220 35 280
rect 55 220 70 280
rect 20 200 70 220
<< ndiffc >>
rect -230 45 -210 105
rect -165 45 -145 105
rect -30 45 -10 105
rect 35 45 55 105
<< pdiffc >>
rect -230 220 -210 280
rect -165 220 -145 280
rect -30 220 -10 280
rect 35 220 55 280
<< psubdiff >>
rect -295 110 -245 125
rect -295 40 -280 110
rect -255 40 -245 110
rect -295 25 -245 40
rect -95 110 -45 125
rect -95 40 -80 110
rect -55 40 -45 110
rect -95 25 -45 40
<< nsubdiff >>
rect -295 285 -245 300
rect -295 215 -280 285
rect -255 215 -245 285
rect -295 200 -245 215
rect -95 285 -45 300
rect -95 215 -80 285
rect -55 215 -45 285
rect -95 200 -45 215
<< psubdiffcont >>
rect -280 40 -255 110
rect -80 40 -55 110
<< nsubdiffcont >>
rect -280 215 -255 285
rect -80 215 -55 285
<< poly >>
rect -195 300 -180 315
rect 5 300 20 315
rect -195 125 -180 200
rect 5 125 20 200
rect -195 10 -180 25
rect 5 10 20 25
rect -220 0 -180 10
rect -220 -20 -210 0
rect -190 -20 -180 0
rect -220 -30 -180 -20
rect -20 0 20 10
rect -20 -20 -10 0
rect 10 -20 20 0
rect -20 -30 20 -20
<< polycont >>
rect -210 -20 -190 0
rect -10 -20 10 0
<< locali >>
rect -290 285 -200 295
rect -290 215 -280 285
rect -255 280 -200 285
rect -255 220 -230 280
rect -210 220 -200 280
rect -255 215 -200 220
rect -290 205 -200 215
rect -175 280 -135 295
rect -175 220 -165 280
rect -145 220 -135 280
rect -175 205 -135 220
rect -90 285 0 295
rect -90 215 -80 285
rect -55 280 0 285
rect -55 220 -30 280
rect -10 220 0 280
rect -55 215 0 220
rect -90 205 0 215
rect 25 280 65 295
rect 25 220 35 280
rect 55 220 65 280
rect 25 205 65 220
rect -160 120 -143 205
rect 40 120 57 205
rect -290 110 -200 120
rect -290 40 -280 110
rect -255 105 -200 110
rect -255 45 -230 105
rect -210 45 -200 105
rect -255 40 -200 45
rect -290 30 -200 40
rect -175 105 -135 120
rect -175 45 -165 105
rect -145 45 -135 105
rect -175 30 -135 45
rect -90 110 0 120
rect -90 40 -80 110
rect -55 105 0 110
rect -55 45 -30 105
rect -10 45 0 105
rect -55 40 0 45
rect -90 30 0 40
rect 25 105 65 120
rect 25 45 35 105
rect 55 45 65 105
rect 25 30 65 45
rect -155 10 -135 30
rect 45 10 65 30
rect -315 0 -180 10
rect -315 -10 -210 0
rect -220 -20 -210 -10
rect -190 -20 -180 0
rect -155 0 20 10
rect -155 -10 -10 0
rect -220 -30 -180 -20
rect -20 -20 -10 -10
rect 10 -20 20 0
rect 45 -10 90 10
rect -20 -30 20 -20
<< viali >>
rect -280 215 -255 285
rect -230 220 -210 280
rect -80 215 -55 285
rect -30 220 -10 280
rect -280 40 -255 110
rect -230 45 -210 105
rect -80 40 -55 110
rect -30 45 -10 105
<< metal1 >>
rect -315 285 90 295
rect -315 215 -280 285
rect -255 280 -80 285
rect -255 220 -230 280
rect -210 220 -80 280
rect -255 215 -80 220
rect -55 280 90 285
rect -55 220 -30 280
rect -10 220 90 280
rect -55 215 90 220
rect -315 205 90 215
rect -315 110 90 120
rect -315 40 -280 110
rect -255 105 -80 110
rect -255 45 -230 105
rect -210 45 -80 105
rect -255 40 -80 45
rect -55 105 90 110
rect -55 45 -30 105
rect -10 45 90 105
rect -55 40 90 45
rect -315 30 90 40
<< labels >>
rlabel metal1 -315 252 -315 252 3 VP
port 3 e
rlabel metal1 -315 47 -315 47 3 VN
port 4 e
rlabel locali -315 0 -315 0 7 A
port 1 w
rlabel locali 90 4 90 4 3 Y
port 2 e
<< end >>
